module sim_cpu
(
      input  wire        clk,
      input  wire        i_rst,
      input  wire        i_timer_irq,

      output wire [31:0] o_ibus_adr,
      output wire        o_ibus_cyc,
      input  wire        i_ibus_gnt,
      input  wire [31:0] i_ibus_rdt,
      input  wire        i_ibus_ack,

      output wire [31:0] o_dbus_adr,
      output wire [31:0] o_dbus_dat,
      output wire        o_dbus_we,
      output wire [3:0]  o_dbus_be,
      output wire        o_dbus_cyc,
      input  wire        i_dbus_gnt,
      input  wire [31:0] i_dbus_rdt,
      input  wire        i_dbus_ack,
      output wire o_core_sleep
//      output wire [31:0] o_debug_req_i,
);

/*   ibex_top cpu
     (.clk_i (clk),
      .rst_ni (!i_rst),

      .test_en_i (1'b1),
      .ram_cfg_i (10'b0),
      .hart_id_i (32'b0),
      .boot_addr_i (32'b0),

      .instr_req_o (o_ibus_cyc),
      .instr_gnt_i (i_ibus_gnt),
      .instr_rvalid_i (i_ibus_ack),
      .instr_addr_o (o_ibus_adr),
      .instr_rdata_i (i_ibus_rdt),
      .instr_rdata_intg_i (7'b0),
      .instr_err_i (1'b0),

      .data_req_o (o_dbus_cyc),
      .data_gnt_i (i_dbus_gnt),
      .data_rvalid_i (i_dbus_ack),
      .data_we_o (o_dbus_we),
      .data_be_o (o_dbus_be), 
      .data_addr_o (o_dbus_adr),
      .data_wdata_o (o_dbus_dat),
      .data_wdata_intg_o (),
      .data_rdata_i (i_dbus_rdt),
      .data_rdata_intg_i (7'b0),
      .data_err_i (1'b0),

      .irq_software_i (1'b0),
      .irq_timer_i (i_timer_irq),
      .irq_external_i (1'b0),
      .irq_fast_i (15'b0),
      .irq_nm_i (1'b0),

      .scramble_key_valid_i (1'b0),
      .scramble_key_i (128'b0),
      .scramble_nonce_i (64'b0),
      .scramble_req_o (),
      .debug_req_i (1'b0),
      .crash_dump_o (),
      .double_fault_seen_o (),
      .fetch_enable_i (4'b0101), // IbexMuBiOn
      .alert_minor_o (),
      .alert_major_internal_o (),
      .alert_major_bus_o (),
      .core_sleep_o (o_core_sleep),
      .scan_rst_ni (1'b1)
   );
*/
  ibex_top cpu (
    .\data_wdata_intg_o[0] (),
    .\data_wdata_intg_o[1] (),
    .\data_wdata_intg_o[2] (),
    .\data_wdata_intg_o[3] (),
    .\data_wdata_intg_o[4] (),
    .\data_wdata_intg_o[5] (),
    .\data_wdata_intg_o[6] (),
    .\scramble_req_o (),
    .\crash_dump_o[0] (),
.\crash_dump_o[1] (),
.\crash_dump_o[2] (),
.\crash_dump_o[3] (),
.\crash_dump_o[4] (),
.\crash_dump_o[5] (),
.\crash_dump_o[6] (),
.\crash_dump_o[7] (),
.\crash_dump_o[8] (),
.\crash_dump_o[9] (),
.\crash_dump_o[10] (),
.\crash_dump_o[11] (),
.\crash_dump_o[12] (),
.\crash_dump_o[13] (),
.\crash_dump_o[14] (),
.\crash_dump_o[15] (),
.\crash_dump_o[16] (),
.\crash_dump_o[17] (),
.\crash_dump_o[18] (),
.\crash_dump_o[19] (),
.\crash_dump_o[20] (),
.\crash_dump_o[21] (),
.\crash_dump_o[22] (),
.\crash_dump_o[23] (),
.\crash_dump_o[24] (),
.\crash_dump_o[25] (),
.\crash_dump_o[26] (),
.\crash_dump_o[27] (),
.\crash_dump_o[28] (),
.\crash_dump_o[29] (),
.\crash_dump_o[30] (),
.\crash_dump_o[31] (),
.\crash_dump_o[32] (),
.\crash_dump_o[33] (),
.\crash_dump_o[34] (),
.\crash_dump_o[35] (),
.\crash_dump_o[36] (),
.\crash_dump_o[37] (),
.\crash_dump_o[38] (),
.\crash_dump_o[39] (),
.\crash_dump_o[40] (),
.\crash_dump_o[41] (),
.\crash_dump_o[42] (),
.\crash_dump_o[43] (),
.\crash_dump_o[44] (),
.\crash_dump_o[45] (),
.\crash_dump_o[46] (),
.\crash_dump_o[47] (),
.\crash_dump_o[48] (),
.\crash_dump_o[49] (),
.\crash_dump_o[50] (),
.\crash_dump_o[51] (),
.\crash_dump_o[52] (),
.\crash_dump_o[53] (),
.\crash_dump_o[54] (),
.\crash_dump_o[55] (),
.\crash_dump_o[56] (),
.\crash_dump_o[57] (),
.\crash_dump_o[58] (),
.\crash_dump_o[59] (),
.\crash_dump_o[60] (),
.\crash_dump_o[61] (),
.\crash_dump_o[62] (),
.\crash_dump_o[63] (),
.\crash_dump_o[64] (),
.\crash_dump_o[65] (),
.\crash_dump_o[66] (),
.\crash_dump_o[67] (),
.\crash_dump_o[68] (),
.\crash_dump_o[69] (),
.\crash_dump_o[70] (),
.\crash_dump_o[71] (),
.\crash_dump_o[72] (),
.\crash_dump_o[73] (),
.\crash_dump_o[74] (),
.\crash_dump_o[75] (),
.\crash_dump_o[76] (),
.\crash_dump_o[77] (),
.\crash_dump_o[78] (),
.\crash_dump_o[79] (),
.\crash_dump_o[80] (),
.\crash_dump_o[81] (),
.\crash_dump_o[82] (),
.\crash_dump_o[83] (),
.\crash_dump_o[84] (),
.\crash_dump_o[85] (),
.\crash_dump_o[86] (),
.\crash_dump_o[87] (),
.\crash_dump_o[88] (),
.\crash_dump_o[89] (),
.\crash_dump_o[90] (),
.\crash_dump_o[91] (),
.\crash_dump_o[92] (),
.\crash_dump_o[93] (),
.\crash_dump_o[94] (),
.\crash_dump_o[95] (),
.\crash_dump_o[96] (),
.\crash_dump_o[97] (),
.\crash_dump_o[98] (),
.\crash_dump_o[99] (),
.\crash_dump_o[100] (),
.\crash_dump_o[101] (),
.\crash_dump_o[102] (),
.\crash_dump_o[103] (),
.\crash_dump_o[104] (),
.\crash_dump_o[105] (),
.\crash_dump_o[106] (),
.\crash_dump_o[107] (),
.\crash_dump_o[108] (),
.\crash_dump_o[109] (),
.\crash_dump_o[110] (),
.\crash_dump_o[111] (),
.\crash_dump_o[112] (),
.\crash_dump_o[113] (),
.\crash_dump_o[114] (),
.\crash_dump_o[115] (),
.\crash_dump_o[116] (),
.\crash_dump_o[117] (),
.\crash_dump_o[118] (),
.\crash_dump_o[119] (),
.\crash_dump_o[120] (),
.\crash_dump_o[121] (),
.\crash_dump_o[122] (),
.\crash_dump_o[123] (),
.\crash_dump_o[124] (),
.\crash_dump_o[125] (),
.\crash_dump_o[126] (),
.\crash_dump_o[127] (),
.\crash_dump_o[128] (),
.\crash_dump_o[129] (),
.\crash_dump_o[130] (),
.\crash_dump_o[131] (),
.\crash_dump_o[132] (),
.\crash_dump_o[133] (),
.\crash_dump_o[134] (),
.\crash_dump_o[135] (),
.\crash_dump_o[136] (),
.\crash_dump_o[137] (),
.\crash_dump_o[138] (),
.\crash_dump_o[139] (),
.\crash_dump_o[140] (),
.\crash_dump_o[141] (),
.\crash_dump_o[142] (),
.\crash_dump_o[143] (),
.\crash_dump_o[144] (),
.\crash_dump_o[145] (),
.\crash_dump_o[146] (),
.\crash_dump_o[147] (),
.\crash_dump_o[148] (),
.\crash_dump_o[149] (),
.\crash_dump_o[150] (),
.\crash_dump_o[151] (),
.\crash_dump_o[152] (),
.\crash_dump_o[153] (),
.\crash_dump_o[154] (),
.\crash_dump_o[155] (),
.\crash_dump_o[156] (),
.\crash_dump_o[157] (),
.\crash_dump_o[158] (),
.\crash_dump_o[159] (),
.\double_fault_seen_o (),
.\alert_minor_o (),
.\alert_major_internal_o (),
.\alert_major_bus_o (),
    .\boot_addr_i[0] (1'h0),
    .\boot_addr_i[10] (1'h0),
    .\boot_addr_i[11] (1'h0),
    .\boot_addr_i[12] (1'h0),
    .\boot_addr_i[13] (1'h0),
    .\boot_addr_i[14] (1'h0),
    .\boot_addr_i[15] (1'h0),
    .\boot_addr_i[16] (1'h0),
    .\boot_addr_i[17] (1'h0),
    .\boot_addr_i[18] (1'h0),
    .\boot_addr_i[19] (1'h0),
    .\boot_addr_i[1] (1'h0),
    .\boot_addr_i[20] (1'h0),
    .\boot_addr_i[21] (1'h0),
    .\boot_addr_i[22] (1'h0),
    .\boot_addr_i[23] (1'h0),
    .\boot_addr_i[24] (1'h0),
    .\boot_addr_i[25] (1'h0),
    .\boot_addr_i[26] (1'h0),
    .\boot_addr_i[27] (1'h0),
    .\boot_addr_i[28] (1'h0),
    .\boot_addr_i[29] (1'h0),
    .\boot_addr_i[2] (1'h0),
    .\boot_addr_i[30] (1'h0),
    .\boot_addr_i[31] (1'h0),
    .\boot_addr_i[3] (1'h0),
    .\boot_addr_i[4] (1'h0),
    .\boot_addr_i[5] (1'h0),
    .\boot_addr_i[6] (1'h0),
    .\boot_addr_i[7] (1'h0),
    .\boot_addr_i[8] (1'h0),
    .\boot_addr_i[9] (1'h0),
    .clk_i(clk),
    .core_sleep_o(o_core_sleep),
    .\data_addr_o[0] (o_dbus_adr[0] ),
    .\data_addr_o[10] (o_dbus_adr[10] ),
    .\data_addr_o[11] (o_dbus_adr[11] ),
    .\data_addr_o[12] (o_dbus_adr[12] ),
    .\data_addr_o[13] (o_dbus_adr[13] ),
    .\data_addr_o[14] (o_dbus_adr[14] ),
    .\data_addr_o[15] (o_dbus_adr[15] ),
    .\data_addr_o[16] (o_dbus_adr[16] ),
    .\data_addr_o[17] (o_dbus_adr[17] ),
    .\data_addr_o[18] (o_dbus_adr[18] ),
    .\data_addr_o[19] (o_dbus_adr[19] ),
    .\data_addr_o[1] (o_dbus_adr[1] ),
    .\data_addr_o[20] (o_dbus_adr[20] ),
    .\data_addr_o[21] (o_dbus_adr[21] ),
    .\data_addr_o[22] (o_dbus_adr[22] ),
    .\data_addr_o[23] (o_dbus_adr[23] ),
    .\data_addr_o[24] (o_dbus_adr[24] ),
    .\data_addr_o[25] (o_dbus_adr[25] ),
    .\data_addr_o[26] (o_dbus_adr[26] ),
    .\data_addr_o[27] (o_dbus_adr[27] ),
    .\data_addr_o[28] (o_dbus_adr[28] ),
    .\data_addr_o[29] (o_dbus_adr[29] ),
    .\data_addr_o[2] (o_dbus_adr[2] ),
    .\data_addr_o[30] (o_dbus_adr[30] ),
    .\data_addr_o[31] (o_dbus_adr[31] ),
    .\data_addr_o[3] (o_dbus_adr[3] ),
    .\data_addr_o[4] (o_dbus_adr[4] ),
    .\data_addr_o[5] (o_dbus_adr[5] ),
    .\data_addr_o[6] (o_dbus_adr[6] ),
    .\data_addr_o[7] (o_dbus_adr[7] ),
    .\data_addr_o[8] (o_dbus_adr[8] ),
    .\data_addr_o[9] (o_dbus_adr[9] ),
    .\data_be_o[0] (o_dbus_be[0] ),
    .\data_be_o[1] (o_dbus_be[1] ),
    .\data_be_o[2] (o_dbus_be[2] ),
    .\data_be_o[3] (o_dbus_be[3] ),
    .data_err_i(1'h0),
    .data_gnt_i(i_dbus_gnt),
    .\data_rdata_i[0] (i_dbus_rdt[0] ),
    .\data_rdata_i[10] (i_dbus_rdt[10] ),
    .\data_rdata_i[11] (i_dbus_rdt[11] ),
    .\data_rdata_i[12] (i_dbus_rdt[12] ),
    .\data_rdata_i[13] (i_dbus_rdt[13] ),
    .\data_rdata_i[14] (i_dbus_rdt[14] ),
    .\data_rdata_i[15] (i_dbus_rdt[15] ),
    .\data_rdata_i[16] (i_dbus_rdt[16] ),
    .\data_rdata_i[17] (i_dbus_rdt[17] ),
    .\data_rdata_i[18] (i_dbus_rdt[18] ),
    .\data_rdata_i[19] (i_dbus_rdt[19] ),
    .\data_rdata_i[1] (i_dbus_rdt[1] ),
    .\data_rdata_i[20] (i_dbus_rdt[20] ),
    .\data_rdata_i[21] (i_dbus_rdt[21] ),
    .\data_rdata_i[22] (i_dbus_rdt[22] ),
    .\data_rdata_i[23] (i_dbus_rdt[23] ),
    .\data_rdata_i[24] (i_dbus_rdt[24] ),
    .\data_rdata_i[25] (i_dbus_rdt[25] ),
    .\data_rdata_i[26] (i_dbus_rdt[26] ),
    .\data_rdata_i[27] (i_dbus_rdt[27] ),
    .\data_rdata_i[28] (i_dbus_rdt[28] ),
    .\data_rdata_i[29] (i_dbus_rdt[29] ),
    .\data_rdata_i[2] (i_dbus_rdt[2] ),
    .\data_rdata_i[30] (i_dbus_rdt[30] ),
    .\data_rdata_i[31] (i_dbus_rdt[31] ),
    .\data_rdata_i[3] (i_dbus_rdt[3] ),
    .\data_rdata_i[4] (i_dbus_rdt[4] ),
    .\data_rdata_i[5] (i_dbus_rdt[5] ),
    .\data_rdata_i[6] (i_dbus_rdt[6] ),
    .\data_rdata_i[7] (i_dbus_rdt[7] ),
    .\data_rdata_i[8] (i_dbus_rdt[8] ),
    .\data_rdata_i[9] (i_dbus_rdt[9] ),
    .\data_rdata_intg_i[0] (1'h0),
    .\data_rdata_intg_i[1] (1'h0),
    .\data_rdata_intg_i[2] (1'h0),
    .\data_rdata_intg_i[3] (1'h0),
    .\data_rdata_intg_i[4] (1'h0),
    .\data_rdata_intg_i[5] (1'h0),
    .\data_rdata_intg_i[6] (1'h0),
    .data_req_o(o_dbus_cyc),
    .data_rvalid_i(i_dbus_ack),
    .\data_wdata_o[0] (o_dbus_dat[0] ),
    .\data_wdata_o[10] (o_dbus_dat[10] ),
    .\data_wdata_o[11] (o_dbus_dat[11] ),
    .\data_wdata_o[12] (o_dbus_dat[12] ),
    .\data_wdata_o[13] (o_dbus_dat[13] ),
    .\data_wdata_o[14] (o_dbus_dat[14] ),
    .\data_wdata_o[15] (o_dbus_dat[15] ),
    .\data_wdata_o[16] (o_dbus_dat[16] ),
    .\data_wdata_o[17] (o_dbus_dat[17] ),
    .\data_wdata_o[18] (o_dbus_dat[18] ),
    .\data_wdata_o[19] (o_dbus_dat[19] ),
    .\data_wdata_o[1] (o_dbus_dat[1] ),
    .\data_wdata_o[20] (o_dbus_dat[20] ),
    .\data_wdata_o[21] (o_dbus_dat[21] ),
    .\data_wdata_o[22] (o_dbus_dat[22] ),
    .\data_wdata_o[23] (o_dbus_dat[23] ),
    .\data_wdata_o[24] (o_dbus_dat[24] ),
    .\data_wdata_o[25] (o_dbus_dat[25] ),
    .\data_wdata_o[26] (o_dbus_dat[26] ),
    .\data_wdata_o[27] (o_dbus_dat[27] ),
    .\data_wdata_o[28] (o_dbus_dat[28] ),
    .\data_wdata_o[29] (o_dbus_dat[29] ),
    .\data_wdata_o[2] (o_dbus_dat[2] ),
    .\data_wdata_o[30] (o_dbus_dat[30] ),
    .\data_wdata_o[31] (o_dbus_dat[31] ),
    .\data_wdata_o[3] (o_dbus_dat[3] ),
    .\data_wdata_o[4] (o_dbus_dat[4] ),
    .\data_wdata_o[5] (o_dbus_dat[5] ),
    .\data_wdata_o[6] (o_dbus_dat[6] ),
    .\data_wdata_o[7] (o_dbus_dat[7] ),
    .\data_wdata_o[8] (o_dbus_dat[8] ),
    .\data_wdata_o[9] (o_dbus_dat[9] ),
    .data_we_o(o_dbus_we),
    .debug_req_i(1'h0),
    .\fetch_enable_i[0] (1'h1),
    .\fetch_enable_i[1] (1'h0),
    .\fetch_enable_i[2] (1'h1),
    .\fetch_enable_i[3] (1'h0),
    .\hart_id_i[0] (1'h0),
    .\hart_id_i[10] (1'h0),
    .\hart_id_i[11] (1'h0),
    .\hart_id_i[12] (1'h0),
    .\hart_id_i[13] (1'h0),
    .\hart_id_i[14] (1'h0),
    .\hart_id_i[15] (1'h0),
    .\hart_id_i[16] (1'h0),
    .\hart_id_i[17] (1'h0),
    .\hart_id_i[18] (1'h0),
    .\hart_id_i[19] (1'h0),
    .\hart_id_i[1] (1'h0),
    .\hart_id_i[20] (1'h0),
    .\hart_id_i[21] (1'h0),
    .\hart_id_i[22] (1'h0),
    .\hart_id_i[23] (1'h0),
    .\hart_id_i[24] (1'h0),
    .\hart_id_i[25] (1'h0),
    .\hart_id_i[26] (1'h0),
    .\hart_id_i[27] (1'h0),
    .\hart_id_i[28] (1'h0),
    .\hart_id_i[29] (1'h0),
    .\hart_id_i[2] (1'h0),
    .\hart_id_i[30] (1'h0),
    .\hart_id_i[31] (1'h0),
    .\hart_id_i[3] (1'h0),
    .\hart_id_i[4] (1'h0),
    .\hart_id_i[5] (1'h0),
    .\hart_id_i[6] (1'h0),
    .\hart_id_i[7] (1'h0),
    .\hart_id_i[8] (1'h0),
    .\hart_id_i[9] (1'h0),
    .\instr_addr_o[0] (o_ibus_adr[0] ),
    .\instr_addr_o[10] (o_ibus_adr[10] ),
    .\instr_addr_o[11] (o_ibus_adr[11] ),
    .\instr_addr_o[12] (o_ibus_adr[12] ),
    .\instr_addr_o[13] (o_ibus_adr[13] ),
    .\instr_addr_o[14] (o_ibus_adr[14] ),
    .\instr_addr_o[15] (o_ibus_adr[15] ),
    .\instr_addr_o[16] (o_ibus_adr[16] ),
    .\instr_addr_o[17] (o_ibus_adr[17] ),
    .\instr_addr_o[18] (o_ibus_adr[18] ),
    .\instr_addr_o[19] (o_ibus_adr[19] ),
    .\instr_addr_o[1] (o_ibus_adr[1] ),
    .\instr_addr_o[20] (o_ibus_adr[20] ),
    .\instr_addr_o[21] (o_ibus_adr[21] ),
    .\instr_addr_o[22] (o_ibus_adr[22] ),
    .\instr_addr_o[23] (o_ibus_adr[23] ),
    .\instr_addr_o[24] (o_ibus_adr[24] ),
    .\instr_addr_o[25] (o_ibus_adr[25] ),
    .\instr_addr_o[26] (o_ibus_adr[26] ),
    .\instr_addr_o[27] (o_ibus_adr[27] ),
    .\instr_addr_o[28] (o_ibus_adr[28] ),
    .\instr_addr_o[29] (o_ibus_adr[29] ),
    .\instr_addr_o[2] (o_ibus_adr[2] ),
    .\instr_addr_o[30] (o_ibus_adr[30] ),
    .\instr_addr_o[31] (o_ibus_adr[31] ),
    .\instr_addr_o[3] (o_ibus_adr[3] ),
    .\instr_addr_o[4] (o_ibus_adr[4] ),
    .\instr_addr_o[5] (o_ibus_adr[5] ),
    .\instr_addr_o[6] (o_ibus_adr[6] ),
    .\instr_addr_o[7] (o_ibus_adr[7] ),
    .\instr_addr_o[8] (o_ibus_adr[8] ),
    .\instr_addr_o[9] (o_ibus_adr[9] ),
    .instr_err_i(1'h0),
    .instr_gnt_i(i_ibus_gnt),
    .\instr_rdata_i[0] (i_ibus_rdt[0] ),
    .\instr_rdata_i[10] (i_ibus_rdt[10] ),
    .\instr_rdata_i[11] (i_ibus_rdt[11] ),
    .\instr_rdata_i[12] (i_ibus_rdt[12] ),
    .\instr_rdata_i[13] (i_ibus_rdt[13] ),
    .\instr_rdata_i[14] (i_ibus_rdt[14] ),
    .\instr_rdata_i[15] (i_ibus_rdt[15] ),
    .\instr_rdata_i[16] (i_ibus_rdt[16] ),
    .\instr_rdata_i[17] (i_ibus_rdt[17] ),
    .\instr_rdata_i[18] (i_ibus_rdt[18] ),
    .\instr_rdata_i[19] (i_ibus_rdt[19] ),
    .\instr_rdata_i[1] (i_ibus_rdt[1] ),
    .\instr_rdata_i[20] (i_ibus_rdt[20] ),
    .\instr_rdata_i[21] (i_ibus_rdt[21] ),
    .\instr_rdata_i[22] (i_ibus_rdt[22] ),
    .\instr_rdata_i[23] (i_ibus_rdt[23] ),
    .\instr_rdata_i[24] (i_ibus_rdt[24] ),
    .\instr_rdata_i[25] (i_ibus_rdt[25] ),
    .\instr_rdata_i[26] (i_ibus_rdt[26] ),
    .\instr_rdata_i[27] (i_ibus_rdt[27] ),
    .\instr_rdata_i[28] (i_ibus_rdt[28] ),
    .\instr_rdata_i[29] (i_ibus_rdt[29] ),
    .\instr_rdata_i[2] (i_ibus_rdt[2] ),
    .\instr_rdata_i[30] (i_ibus_rdt[30] ),
    .\instr_rdata_i[31] (i_ibus_rdt[31] ),
    .\instr_rdata_i[3] (i_ibus_rdt[3] ),
    .\instr_rdata_i[4] (i_ibus_rdt[4] ),
    .\instr_rdata_i[5] (i_ibus_rdt[5] ),
    .\instr_rdata_i[6] (i_ibus_rdt[6] ),
    .\instr_rdata_i[7] (i_ibus_rdt[7] ),
    .\instr_rdata_i[8] (i_ibus_rdt[8] ),
    .\instr_rdata_i[9] (i_ibus_rdt[9] ),
    .\instr_rdata_intg_i[0] (1'h0),
    .\instr_rdata_intg_i[1] (1'h0),
    .\instr_rdata_intg_i[2] (1'h0),
    .\instr_rdata_intg_i[3] (1'h0),
    .\instr_rdata_intg_i[4] (1'h0),
    .\instr_rdata_intg_i[5] (1'h0),
    .\instr_rdata_intg_i[6] (1'h0),
    .instr_req_o(o_ibus_cyc),
    .instr_rvalid_i(i_ibus_ack),
    .irq_external_i(1'h0),
    .\irq_fast_i[0] (1'h0),
    .\irq_fast_i[10] (1'h0),
    .\irq_fast_i[11] (1'h0),
    .\irq_fast_i[12] (1'h0),
    .\irq_fast_i[13] (1'h0),
    .\irq_fast_i[14] (1'h0),
    .\irq_fast_i[1] (1'h0),
    .\irq_fast_i[2] (1'h0),
    .\irq_fast_i[3] (1'h0),
    .\irq_fast_i[4] (1'h0),
    .\irq_fast_i[5] (1'h0),
    .\irq_fast_i[6] (1'h0),
    .\irq_fast_i[7] (1'h0),
    .\irq_fast_i[8] (1'h0),
    .\irq_fast_i[9] (1'h0),
    .irq_nm_i(1'h0),
    .irq_software_i(1'h0),
    .irq_timer_i(i_timer_irq),
    .\ram_cfg_i[0] (1'h0),
    .\ram_cfg_i[1] (1'h0),
    .\ram_cfg_i[2] (1'h0),
    .\ram_cfg_i[3] (1'h0),
    .\ram_cfg_i[4] (1'h0),
    .\ram_cfg_i[5] (1'h0),
    .\ram_cfg_i[6] (1'h0),
    .\ram_cfg_i[7] (1'h0),
    .\ram_cfg_i[8] (1'h0),
    .\ram_cfg_i[9] (1'h0),
    .rst_ni (!i_rst),
    .scan_rst_ni(1'h1),
    .\scramble_key_i[0] (1'h0),
    .\scramble_key_i[100] (1'h0),
    .\scramble_key_i[101] (1'h0),
    .\scramble_key_i[102] (1'h0),
    .\scramble_key_i[103] (1'h0),
    .\scramble_key_i[104] (1'h0),
    .\scramble_key_i[105] (1'h0),
    .\scramble_key_i[106] (1'h0),
    .\scramble_key_i[107] (1'h0),
    .\scramble_key_i[108] (1'h0),
    .\scramble_key_i[109] (1'h0),
    .\scramble_key_i[10] (1'h0),
    .\scramble_key_i[110] (1'h0),
    .\scramble_key_i[111] (1'h0),
    .\scramble_key_i[112] (1'h0),
    .\scramble_key_i[113] (1'h0),
    .\scramble_key_i[114] (1'h0),
    .\scramble_key_i[115] (1'h0),
    .\scramble_key_i[116] (1'h0),
    .\scramble_key_i[117] (1'h0),
    .\scramble_key_i[118] (1'h0),
    .\scramble_key_i[119] (1'h0),
    .\scramble_key_i[11] (1'h0),
    .\scramble_key_i[120] (1'h0),
    .\scramble_key_i[121] (1'h0),
    .\scramble_key_i[122] (1'h0),
    .\scramble_key_i[123] (1'h0),
    .\scramble_key_i[124] (1'h0),
    .\scramble_key_i[125] (1'h0),
    .\scramble_key_i[126] (1'h0),
    .\scramble_key_i[127] (1'h0),
    .\scramble_key_i[12] (1'h0),
    .\scramble_key_i[13] (1'h0),
    .\scramble_key_i[14] (1'h0),
    .\scramble_key_i[15] (1'h0),
    .\scramble_key_i[16] (1'h0),
    .\scramble_key_i[17] (1'h0),
    .\scramble_key_i[18] (1'h0),
    .\scramble_key_i[19] (1'h0),
    .\scramble_key_i[1] (1'h0),
    .\scramble_key_i[20] (1'h0),
    .\scramble_key_i[21] (1'h0),
    .\scramble_key_i[22] (1'h0),
    .\scramble_key_i[23] (1'h0),
    .\scramble_key_i[24] (1'h0),
    .\scramble_key_i[25] (1'h0),
    .\scramble_key_i[26] (1'h0),
    .\scramble_key_i[27] (1'h0),
    .\scramble_key_i[28] (1'h0),
    .\scramble_key_i[29] (1'h0),
    .\scramble_key_i[2] (1'h0),
    .\scramble_key_i[30] (1'h0),
    .\scramble_key_i[31] (1'h0),
    .\scramble_key_i[32] (1'h0),
    .\scramble_key_i[33] (1'h0),
    .\scramble_key_i[34] (1'h0),
    .\scramble_key_i[35] (1'h0),
    .\scramble_key_i[36] (1'h0),
    .\scramble_key_i[37] (1'h0),
    .\scramble_key_i[38] (1'h0),
    .\scramble_key_i[39] (1'h0),
    .\scramble_key_i[3] (1'h0),
    .\scramble_key_i[40] (1'h0),
    .\scramble_key_i[41] (1'h0),
    .\scramble_key_i[42] (1'h0),
    .\scramble_key_i[43] (1'h0),
    .\scramble_key_i[44] (1'h0),
    .\scramble_key_i[45] (1'h0),
    .\scramble_key_i[46] (1'h0),
    .\scramble_key_i[47] (1'h0),
    .\scramble_key_i[48] (1'h0),
    .\scramble_key_i[49] (1'h0),
    .\scramble_key_i[4] (1'h0),
    .\scramble_key_i[50] (1'h0),
    .\scramble_key_i[51] (1'h0),
    .\scramble_key_i[52] (1'h0),
    .\scramble_key_i[53] (1'h0),
    .\scramble_key_i[54] (1'h0),
    .\scramble_key_i[55] (1'h0),
    .\scramble_key_i[56] (1'h0),
    .\scramble_key_i[57] (1'h0),
    .\scramble_key_i[58] (1'h0),
    .\scramble_key_i[59] (1'h0),
    .\scramble_key_i[5] (1'h0),
    .\scramble_key_i[60] (1'h0),
    .\scramble_key_i[61] (1'h0),
    .\scramble_key_i[62] (1'h0),
    .\scramble_key_i[63] (1'h0),
    .\scramble_key_i[64] (1'h0),
    .\scramble_key_i[65] (1'h0),
    .\scramble_key_i[66] (1'h0),
    .\scramble_key_i[67] (1'h0),
    .\scramble_key_i[68] (1'h0),
    .\scramble_key_i[69] (1'h0),
    .\scramble_key_i[6] (1'h0),
    .\scramble_key_i[70] (1'h0),
    .\scramble_key_i[71] (1'h0),
    .\scramble_key_i[72] (1'h0),
    .\scramble_key_i[73] (1'h0),
    .\scramble_key_i[74] (1'h0),
    .\scramble_key_i[75] (1'h0),
    .\scramble_key_i[76] (1'h0),
    .\scramble_key_i[77] (1'h0),
    .\scramble_key_i[78] (1'h0),
    .\scramble_key_i[79] (1'h0),
    .\scramble_key_i[7] (1'h0),
    .\scramble_key_i[80] (1'h0),
    .\scramble_key_i[81] (1'h0),
    .\scramble_key_i[82] (1'h0),
    .\scramble_key_i[83] (1'h0),
    .\scramble_key_i[84] (1'h0),
    .\scramble_key_i[85] (1'h0),
    .\scramble_key_i[86] (1'h0),
    .\scramble_key_i[87] (1'h0),
    .\scramble_key_i[88] (1'h0),
    .\scramble_key_i[89] (1'h0),
    .\scramble_key_i[8] (1'h0),
    .\scramble_key_i[90] (1'h0),
    .\scramble_key_i[91] (1'h0),
    .\scramble_key_i[92] (1'h0),
    .\scramble_key_i[93] (1'h0),
    .\scramble_key_i[94] (1'h0),
    .\scramble_key_i[95] (1'h0),
    .\scramble_key_i[96] (1'h0),
    .\scramble_key_i[97] (1'h0),
    .\scramble_key_i[98] (1'h0),
    .\scramble_key_i[99] (1'h0),
    .\scramble_key_i[9] (1'h0),
    .scramble_key_valid_i(1'h0),
    .\scramble_nonce_i[0] (1'h0),
    .\scramble_nonce_i[10] (1'h0),
    .\scramble_nonce_i[11] (1'h0),
    .\scramble_nonce_i[12] (1'h0),
    .\scramble_nonce_i[13] (1'h0),
    .\scramble_nonce_i[14] (1'h0),
    .\scramble_nonce_i[15] (1'h0),
    .\scramble_nonce_i[16] (1'h0),
    .\scramble_nonce_i[17] (1'h0),
    .\scramble_nonce_i[18] (1'h0),
    .\scramble_nonce_i[19] (1'h0),
    .\scramble_nonce_i[1] (1'h0),
    .\scramble_nonce_i[20] (1'h0),
    .\scramble_nonce_i[21] (1'h0),
    .\scramble_nonce_i[22] (1'h0),
    .\scramble_nonce_i[23] (1'h0),
    .\scramble_nonce_i[24] (1'h0),
    .\scramble_nonce_i[25] (1'h0),
    .\scramble_nonce_i[26] (1'h0),
    .\scramble_nonce_i[27] (1'h0),
    .\scramble_nonce_i[28] (1'h0),
    .\scramble_nonce_i[29] (1'h0),
    .\scramble_nonce_i[2] (1'h0),
    .\scramble_nonce_i[30] (1'h0),
    .\scramble_nonce_i[31] (1'h0),
    .\scramble_nonce_i[32] (1'h0),
    .\scramble_nonce_i[33] (1'h0),
    .\scramble_nonce_i[34] (1'h0),
    .\scramble_nonce_i[35] (1'h0),
    .\scramble_nonce_i[36] (1'h0),
    .\scramble_nonce_i[37] (1'h0),
    .\scramble_nonce_i[38] (1'h0),
    .\scramble_nonce_i[39] (1'h0),
    .\scramble_nonce_i[3] (1'h0),
    .\scramble_nonce_i[40] (1'h0),
    .\scramble_nonce_i[41] (1'h0),
    .\scramble_nonce_i[42] (1'h0),
    .\scramble_nonce_i[43] (1'h0),
    .\scramble_nonce_i[44] (1'h0),
    .\scramble_nonce_i[45] (1'h0),
    .\scramble_nonce_i[46] (1'h0),
    .\scramble_nonce_i[47] (1'h0),
    .\scramble_nonce_i[48] (1'h0),
    .\scramble_nonce_i[49] (1'h0),
    .\scramble_nonce_i[4] (1'h0),
    .\scramble_nonce_i[50] (1'h0),
    .\scramble_nonce_i[51] (1'h0),
    .\scramble_nonce_i[52] (1'h0),
    .\scramble_nonce_i[53] (1'h0),
    .\scramble_nonce_i[54] (1'h0),
    .\scramble_nonce_i[55] (1'h0),
    .\scramble_nonce_i[56] (1'h0),
    .\scramble_nonce_i[57] (1'h0),
    .\scramble_nonce_i[58] (1'h0),
    .\scramble_nonce_i[59] (1'h0),
    .\scramble_nonce_i[5] (1'h0),
    .\scramble_nonce_i[60] (1'h0),
    .\scramble_nonce_i[61] (1'h0),
    .\scramble_nonce_i[62] (1'h0),
    .\scramble_nonce_i[63] (1'h0),
    .\scramble_nonce_i[6] (1'h0),
    .\scramble_nonce_i[7] (1'h0),
    .\scramble_nonce_i[8] (1'h0),
    .\scramble_nonce_i[9] (1'h0),
    .test_en_i(1'h1)
  );

endmodule
/*
module ibex_top(
  // Clock and Reset input  logic                         clk_i,
  input  logic                         rst_ni,

  input  logic                         test_en_i,     // enable all clock gates for testing
  input  logic [9:0]  ram_cfg_i,

  input  logic [31:0]                  hart_id_i,
  input  logic [31:0]                  boot_addr_i,

  // Instruction memory interface
  output logic                         instr_req_o,
  input  logic                         instr_gnt_i,
  input  logic                         instr_rvalid_i,
  output logic [31:0]                  instr_addr_o,
  input  logic [31:0]                  instr_rdata_i,
  input  logic [6:0]                   instr_rdata_intg_i,
  input  logic                         instr_err_i,

  // Data memory interface
  output logic                         data_req_o,
  input  logic                         data_gnt_i,
  input  logic                         data_rvalid_i,
  output logic                         data_we_o,
  output logic [3:0]                   data_be_o,
  output logic [31:0]                  data_addr_o,
  output logic [31:0]                  data_wdata_o,
  output logic [6:0]                   data_wdata_intg_o,
  input  logic [31:0]                  data_rdata_i,
  input  logic [6:0]                   data_rdata_intg_i,
  input  logic                         data_err_i,

  // Interrupt inputs
  input  logic                         irq_software_i,
  input  logic                         irq_timer_i,
  input  logic                         irq_external_i,
  input  logic [14:0]                  irq_fast_i,
  input  logic                         irq_nm_i,       // non-maskeable interrupt

  // Scrambling Interface
  input  logic                         scramble_key_valid_i,
  input  logic [128-1:0]    scramble_key_i,
  input  logic [64-1:0]  scramble_nonce_i,
  output logic                         scramble_req_o,

  // Debug Interface
  input  logic                         debug_req_i,
  output logic [159:0]                  crash_dump_o,
  output logic                         double_fault_seen_o,

  // RISC-V Formal Interface
  // Does not comply with the coding standards of _i/_o suffixes, but follows
  // the convention of RISC-V Formal Interface Specification.
`ifdef RVFI
  output logic                         rvfi_valid,
  output logic [63:0]                  rvfi_order,
  output logic [31:0]                  rvfi_insn,
  output logic                         rvfi_trap,
  output logic                         rvfi_halt,
  output logic                         rvfi_intr,
  output logic [ 1:0]                  rvfi_mode,
  output logic [ 1:0]                  rvfi_ixl,
  output logic [ 4:0]                  rvfi_rs1_addr,
  output logic [ 4:0]                  rvfi_rs2_addr,
  output logic [ 4:0]                  rvfi_rs3_addr,
  output logic [31:0]                  rvfi_rs1_rdata,
  output logic [31:0]                  rvfi_rs2_rdata,
  output logic [31:0]                  rvfi_rs3_rdata,
  output logic [ 4:0]                  rvfi_rd_addr,
  output logic [31:0]                  rvfi_rd_wdata,
  output logic [31:0]                  rvfi_pc_rdata,
  output logic [31:0]                  rvfi_pc_wdata,
  output logic [31:0]                  rvfi_mem_addr,
  output logic [ 3:0]                  rvfi_mem_rmask,
  output logic [ 3:0]                  rvfi_mem_wmask,
  output logic [31:0]                  rvfi_mem_rdata,
  output logic [31:0]                  rvfi_mem_wdata,
  output logic [31:0]                  rvfi_ext_mip,
  output logic                         rvfi_ext_nmi,
  output logic                         rvfi_ext_nmi_int,
  output logic                         rvfi_ext_debug_req,
  output logic                         rvfi_ext_debug_mode,
  output logic                         rvfi_ext_rf_wr_suppress,
  output logic [63:0]                  rvfi_ext_mcycle,
  output logic [31:0]                  rvfi_ext_mhpmcounters [10],
  output logic [31:0]                  rvfi_ext_mhpmcountersh [10],
  output logic                         rvfi_ext_ic_scr_key_valid,
  output logic                         rvfi_ext_irq_valid,
`endif

  // CPU Control Signals
  input  logic [3:0]                   fetch_enable_i,
  output logic                         alert_minor_o,
  output logic                         alert_major_internal_o,
  output logic                         alert_major_bus_o,
  output logic                         core_sleep_o,

  // DFT bypass controls
  input logic                          scan_rst_ni
);*/
